/*
############################################# 
# ECE 540 project 2
#
# Author:	Rafael Schultz (srafael@pdx.edu)
# Date:		12-Nov-2023	
#
# Changes made to include VGA peripheral
#
# Targeted to Nexys A7 FPGA board
#############################################
*/



module char_to_pix (
	input wire [7:0]	char_data,
	input wire [3:0]	index,
	output reg [0:15]	pixel_line // 16 bit for the character selected line
);


  // when data or line requested changes, convert to line with 16 pixels
  always @(*) begin 
	case ({char_data, index}) // use the 8 bits of the ASCII character, 4 bits of index because 16 lines
		12'h300: 	pixel_line =  	16'b0001111111100000;  // 0 in ASCII
		12'h301:	pixel_line =  	16'b0011111111110000;
		12'h302:	pixel_line =	16'b0111100001111000;
		12'h303:	pixel_line =	16'b1111000000111100;
		12'h304:	pixel_line =	16'b1111000001111100;
		12'h305:	pixel_line =	16'b1111000011111100;
		12'h306:	pixel_line =	16'b1111000111111100;
		12'h307:	pixel_line =	16'b1111001110111100;
		12'h308:	pixel_line =	16'b1111011100111100;
		12'h309:	pixel_line =	16'b1111111000111100;
		12'h30A:	pixel_line =	16'b1111110000111100;
		12'h30B:	pixel_line =	16'b0111110000111100;
		12'h30C:	pixel_line =	16'b0011111111111000;
		12'h30D:	pixel_line =	16'b0001111111110000;
		12'h30E:	pixel_line =	16'b0000000000000000;
		12'h30F:	pixel_line =	16'b0000000000000000;
		
		12'h310: 	pixel_line =  	16'b0000011100000000;  // 1 in ASCII
		12'h311:	pixel_line =  	16'b0000111100000000;
		12'h312:	pixel_line =	16'b0011111100000000;
		12'h313:	pixel_line =	16'b0111111100000000;
		12'h314:	pixel_line =	16'b0000111100000000;
		12'h315:	pixel_line =	16'b0000111100000000;
		12'h316:	pixel_line =	16'b0000111100000000;
		12'h317:	pixel_line =	16'b0000111100000000;
		12'h318:	pixel_line =	16'b0000111100000000;
		12'h319:	pixel_line =	16'b0000111100000000;
		12'h31A:	pixel_line =	16'b0000111100000000;
		12'h31B:	pixel_line =	16'b0000111100000000;
		12'h31C:	pixel_line =	16'b1111111111110000;
		12'h31D:	pixel_line =	16'b1111111111110000;
		12'h31E:	pixel_line =	16'b0000000000000000;
		12'h31F:	pixel_line =	16'b0000000000000000;
		

		12'h320: 	pixel_line =  	16'b0001111111000000;  // 2 in ASCII
		12'h321:	pixel_line =  	16'b0011111111100000;
		12'h322:	pixel_line =	16'b0111000011110000;
		12'h323:	pixel_line =	16'b1110000011110000;
		12'h324:	pixel_line =	16'b0000000111100000;
		12'h325:	pixel_line =	16'b0000001111000000;
		12'h326:	pixel_line =	16'b0000011110000000;
		12'h327:	pixel_line =	16'b0000111100000000;
		12'h328:	pixel_line =	16'b0001111000000000;
		12'h329:	pixel_line =	16'b0011110000000000;
		12'h32A:	pixel_line =	16'b0111100001110000;
		12'h32B:	pixel_line =	16'b1111000001110000;
		12'h32C:	pixel_line =	16'b1111111111110000;
		12'h32D:	pixel_line =	16'b1111111111110000;
		12'h32E:	pixel_line =	16'b0000000000000000;
		12'h32F:	pixel_line =	16'b0000000000000000;

		12'h330:	pixel_line =  	16'b0001111110000000;  // 3 in ASCII
		12'h331:	pixel_line =  	16'b0011111111000000;
		12'h332:	pixel_line =	16'b0111000111100000;
		12'h333:	pixel_line =	16'b1110000011110000;
		12'h334:	pixel_line =	16'b0000000011110000;
		12'h335:	pixel_line =	16'b0000000111100000;
		12'h336:	pixel_line =	16'b0000111111000000;
		12'h337:	pixel_line =	16'b0000111111000000;
		12'h338:	pixel_line =	16'b0000000111100000;
		12'h339:	pixel_line =	16'b0000000011110000;
		12'h33A:	pixel_line =	16'b1110000011110000;
		12'h33B:	pixel_line =	16'b0111000111100000;
		12'h33C:	pixel_line =	16'b0011111111000000;
		12'h33D:	pixel_line =	16'b0001111110000000;
		12'h33E:	pixel_line =	16'b0000000000000000;
		12'h33F:	pixel_line =	16'b0000000000000000;

		12'h340: 	pixel_line =  	16'b0000000111110000;  // 4 in ASCII	
		12'h341:	pixel_line =  	16'b0000001111110000;
		12'h342:	pixel_line =	16'b0000011111110000;
		12'h343:	pixel_line =	16'b0000111011110000;
		12'h344:	pixel_line =	16'b0001110011110000;
		12'h345:	pixel_line =	16'b0011100011110000;
		12'h346:	pixel_line =	16'b0111000011110000;
		12'h347:	pixel_line =	16'b1110000011110000;
		12'h348:	pixel_line =	16'b1111111111111100;
		12'h349:	pixel_line =	16'b1111111111111100;
		12'h34A:	pixel_line =	16'b0000000011110000;
		12'h34B:	pixel_line =	16'b0000000011110000;
		12'h34C:	pixel_line =	16'b0000001111111100;
		12'h34D:	pixel_line =	16'b0000001111111100;
		12'h34E:	pixel_line =	16'b0000000000000000;
		12'h34F:	pixel_line =	16'b0000000000000000;

		12'h350: 	pixel_line =  	16'b1111111111110000;  // 5 in ASCII
		12'h351:	pixel_line =  	16'b1111111111110000;
		12'h352:	pixel_line =	16'b1111000000000000;
		12'h353:	pixel_line =	16'b1111000000000000;
		12'h354:	pixel_line =	16'b1111111110000000;
		12'h355:	pixel_line =	16'b1111111111000000;
		12'h356:	pixel_line =	16'b0000000111110000;
		12'h357:	pixel_line =	16'b0000000011110000;
		12'h358:	pixel_line =	16'b0000000011110000;
		12'h359:	pixel_line =	16'b0000000011110000;
		12'h35A:	pixel_line =	16'b1110000011110000;
		12'h35B:	pixel_line =	16'b1111000011110000;
		12'h35C:	pixel_line =	16'b0111111111100000;
		12'h35D:	pixel_line =	16'b0011111111000000;
		12'h35E:	pixel_line =	16'b0000000000000000;
		12'h35F:	pixel_line =	16'b0000000000000000;

		12'h360: 	pixel_line =  	16'b0000011111000000;  // 6 in ASCII
		12'h361:	pixel_line =  	16'b0000111111000000;
		12'h362:	pixel_line =	16'b0011111000000000;
		12'h363:	pixel_line =	16'b0011110000000000;
		12'h364:	pixel_line =	16'b0111100000000000;
		12'h365:	pixel_line =	16'b1111000000000000;
		12'h366:	pixel_line =	16'b1111111100000000;
		12'h367:	pixel_line =	16'b1111111111000000;
		12'h368:	pixel_line =	16'b1111000011110000;
		12'h369:	pixel_line =	16'b1111000011110000;
		12'h36A:	pixel_line =	16'b1111000011110000;
		12'h36B:	pixel_line =	16'b1111000011110000;
		12'h36C:	pixel_line =	16'b0111111111100000;
		12'h36D:	pixel_line =	16'b0011111111000000;
		12'h36E:	pixel_line =	16'b0000000000000000;
		12'h36F:	pixel_line =	16'b0000000000000000;

		12'h370: 	pixel_line =  	16'b1111111111100000;  // 7 in ASCII
		12'h371:	pixel_line =  	16'b1111111111110000;
		12'h372:	pixel_line =	16'b1111000011110000;
		12'h373:	pixel_line =	16'b1111000011110000;
		12'h374:	pixel_line =	16'b0000000011110000;
		12'h375:	pixel_line =	16'b0000000111110000;
		12'h376:	pixel_line =	16'b0000001111100000;
		12'h377:	pixel_line =	16'b0000011111000000;
		12'h378:	pixel_line =	16'b0000111110000000;
		12'h379:	pixel_line =	16'b0000111100000000;
		12'h37A:	pixel_line =	16'b0000111100000000;
		12'h37B:	pixel_line =	16'b0000111100000000;
		12'h37C:	pixel_line =	16'b0000111100000000;
		12'h37D:	pixel_line =	16'b0000111100000000;
		12'h37E:	pixel_line =	16'b0000000000000000;
		12'h37F:	pixel_line =	16'b0000000000000000;

		12'h380: 	pixel_line =  	16'b0001111110000000;  // 8 in ASCII
		12'h381:	pixel_line =  	16'b0111111111100000;
		12'h382:	pixel_line =	16'b1111000011110000;
		12'h383:	pixel_line =	16'b1111000011110000;
		12'h384:	pixel_line =	16'b1111000011110000;
		12'h385:	pixel_line =	16'b0111000011100000;
		12'h386:	pixel_line =	16'b0011111111000000;
		12'h387:	pixel_line =	16'b0011111111000000;
		12'h388:	pixel_line =	16'b0111000011100000;
		12'h389:	pixel_line =	16'b1111000011110000;
		12'h38A:	pixel_line =	16'b1111000011110000;
		12'h38B:	pixel_line =	16'b1111000011110000;
		12'h38C:	pixel_line =	16'b0111111111100000;
		12'h38D:	pixel_line =	16'b0011111111000000;
		12'h38E:	pixel_line =	16'b0000000000000000;
		12'h38F:	pixel_line =	16'b0000000000000000;

		12'h390: 	pixel_line =  	16'b0001111110000000;  // 9 in ASCII	
		12'h391:	pixel_line =  	16'b0011111111000000;
		12'h392:	pixel_line =	16'b0111000011100000;
		12'h393:	pixel_line =	16'b1111000011110000;
		12'h394:	pixel_line =	16'b1111000011110000;
		12'h395:	pixel_line =	16'b1111000011110000;
		12'h396:	pixel_line =	16'b0111111111110000;
		12'h397:	pixel_line =	16'b0011111111110000;
		12'h398:	pixel_line =	16'b0000000111110000;
		12'h399:	pixel_line =	16'b0000000011100000;
		12'h39A:	pixel_line =	16'b0000000111000000;
		12'h39B:	pixel_line =	16'b0000001110000000;
		12'h39C:	pixel_line =	16'b0011111100000000;
		12'h39D:	pixel_line =	16'b0011111000000000;
		12'h39E:	pixel_line =	16'b0000000000000000;
		12'h39F:	pixel_line =	16'b0000000000000000;

		12'h610:	pixel_line =  	16'b0000000000000000;  // a in ASCII
		12'h611:	pixel_line =  	16'b0000000000000000;
		12'h612:	pixel_line =  	16'b0000000000000000;
		12'h613:	pixel_line =  	16'b0000001111100000;
		12'h614:	pixel_line =  	16'b0000111111111000;
		12'h615:	pixel_line =  	16'b0001110001111000;
		12'h616:	pixel_line =  	16'b0011100001110000;
		12'h617:	pixel_line =  	16'b0011100001110000;
		12'h618:	pixel_line =  	16'b0011100001110000;
		12'h619:	pixel_line =  	16'b0011100001110000;
		12'h61A:	pixel_line =  	16'b0011110001111000;
		12'h61B:	pixel_line =  	16'b0001111111011000;
		12'h61C:	pixel_line =  	16'b0000111110011100;
		12'h61D:	pixel_line =  	16'b0000000000000000;
		12'h61E:	pixel_line =  	16'b0000000000000000;
		12'h61F:	pixel_line =  	16'b0000000000000000;


		12'h620:	pixel_line =  	16'b0000000000000000;  // b in ASCII
		12'h621:	pixel_line =  	16'b0011100000000000;
		12'h622:	pixel_line =  	16'b0011100000000000;
		12'h623:	pixel_line =  	16'b0011100110000000;
		12'h624:	pixel_line =  	16'b0011101111100000;
		12'h625:	pixel_line =  	16'b0011111111111000;
		12'h626:	pixel_line =  	16'b0011100000111100;
		12'h627:	pixel_line =  	16'b0011100000011100;
		12'h628:	pixel_line =  	16'b0011100000011100;
		12'h629:	pixel_line =  	16'b0011100000111100;
		12'h62A:	pixel_line =  	16'b0011111111111000;
		12'h62B:	pixel_line =  	16'b0011011111110000;
		12'h62C:	pixel_line =  	16'b0011001111100000;
		12'h62D:	pixel_line =  	16'b0000000000000000;
		12'h62E:	pixel_line =  	16'b0000000000000000;
		12'h62F:	pixel_line =  	16'b0000000000000000;

		12'h630:	pixel_line =  	16'b0000000000000000;  // c in ASCII
		12'h631:	pixel_line =  	16'b0000000000000000;
		12'h632:	pixel_line =  	16'b0000000000000000;
		12'h633:	pixel_line =  	16'b0000011111000000;
		12'h634:	pixel_line =  	16'b0001111111110000;
		12'h635:	pixel_line =  	16'b0011110001111000;
		12'h636:	pixel_line =  	16'b0011110000111000;
		12'h637:	pixel_line =  	16'b0011110000000000;
		12'h638:	pixel_line =  	16'b0011110000000000;
		12'h639:	pixel_line =  	16'b0011110000111000;
		12'h63A:	pixel_line =  	16'b0011110001111000;
		12'h63B:	pixel_line =  	16'b0001111111110000;
		12'h63C:	pixel_line =  	16'b0000111111100000;
		12'h63D:	pixel_line =  	16'b0000000000000000;
		12'h63E:	pixel_line =  	16'b0000000000000000;
		12'h63F:	pixel_line =  	16'b0000000000000000;

		12'h640:	pixel_line =  	16'b0000000000000000;  // d in ASCII
		12'h641:	pixel_line =  	16'b0000000000011100;
		12'h642:	pixel_line =  	16'b0000000000011100;
		12'h643:	pixel_line =  	16'b0000000110011100;
		12'h644:	pixel_line =  	16'b0000111111111100;
		12'h645:	pixel_line =  	16'b0001111111111100;
		12'h646:	pixel_line =  	16'b0011110000011100;
		12'h647:	pixel_line =  	16'b0011100000011100;
		12'h648:	pixel_line =  	16'b0011100000011100;
		12'h649:	pixel_line =  	16'b0011110000011100;
		12'h64A:	pixel_line =  	16'b0001111111111100;
		12'h64B:	pixel_line =  	16'b0000111111101100;
		12'h64C:	pixel_line =  	16'b0000011111001100;
		12'h64D:	pixel_line =  	16'b0000000000000000;
		12'h64E:	pixel_line =  	16'b0000000000000000;
		12'h64F:	pixel_line =  	16'b0000000000000000;

		12'h650:	pixel_line =  	16'b0000000000000000;  // e in ASCII
		12'h651:	pixel_line =  	16'b0000000000000000;
		12'h652:	pixel_line =  	16'b0000000000000000;
		12'h653:	pixel_line =  	16'b0000111111100000;
		12'h654:	pixel_line =  	16'b0001111111110000;
		12'h655:	pixel_line =  	16'b0011110001111000;
		12'h656:	pixel_line =  	16'b0011100000111000;
		12'h657:	pixel_line =  	16'b0011111111110000;
		12'h658:	pixel_line =  	16'b0011110000000000;
		12'h659:	pixel_line =  	16'b0011100000000000;
		12'h65A:	pixel_line =  	16'b0011110000111000;
		12'h65B:	pixel_line =  	16'b0001111111111000;
		12'h65C:	pixel_line =  	16'b0000111111100000;
		12'h65D:	pixel_line =  	16'b0000000000000000;
		12'h65E:	pixel_line =  	16'b0000000000000000;
		12'h65F:	pixel_line =  	16'b0000000000000000;

		12'h660:	pixel_line =  	16'b0000000000000000;  // f in ASCII
		12'h661:	pixel_line =  	16'b0000000111111000;
		12'h662:	pixel_line =  	16'b0000011111111000;
		12'h663:	pixel_line =  	16'b0000111111000000;
		12'h664:	pixel_line =  	16'b0000111100000000;
		12'h665:	pixel_line =  	16'b0000111100000000;
		12'h666:	pixel_line =  	16'b0111111111111000;
		12'h667:	pixel_line =  	16'b0111111111111000;
		12'h668:	pixel_line =  	16'b0000111100000000;
		12'h669:	pixel_line =  	16'b0000111100000000;
		12'h66A:	pixel_line =  	16'b0000111100000000;
		12'h66B:	pixel_line =  	16'b0000111100000000;
		12'h66C:	pixel_line =  	16'b0000111100000000;
		12'h66D:	pixel_line =  	16'b0000111100000000;
		12'h66E:	pixel_line =  	16'b0000000000000000;
		12'h66F:	pixel_line =  	16'b0000000000000000;

		12'h670:	pixel_line =  	16'b0000000000000000;  // g in ASCII
		12'h671:	pixel_line =  	16'b0000000000000000;
		12'h672:	pixel_line =  	16'b0000000000000000;
		12'h673:	pixel_line =  	16'b0000111111111100;
		12'h674:	pixel_line =  	16'b0001110000111000;
		12'h675:	pixel_line =  	16'b0011100000011100;
		12'h676:	pixel_line =  	16'b0011110000111000;
		12'h677:	pixel_line =  	16'b0011111111110000;
		12'h678:	pixel_line =  	16'b0001110000000000;
		12'h679:	pixel_line =  	16'b0001110000000000;
		12'h67A:	pixel_line =  	16'b0001111111110000;
		12'h67B:	pixel_line =  	16'b0011111001111000;
		12'h67C:	pixel_line =  	16'b0011100000111000;
		12'h67D:	pixel_line =  	16'b0001111001111000;
		12'h67E:	pixel_line =  	16'b0000111111100000;
		12'h67F:	pixel_line =  	16'b0000000000000000;

		12'h680:	pixel_line =  	16'b0000000000000000;  // h in ASCII 
		12'h681:	pixel_line =  	16'b0011100000000000;
		12'h682:	pixel_line =  	16'b0011100000000000;
		12'h683:	pixel_line =  	16'b0011100000000000;
		12'h684:	pixel_line =  	16'b0011100000000000;
		12'h685:	pixel_line =  	16'b0011101100000000;
		12'h686:	pixel_line =  	16'b0011111111000000;
		12'h687:	pixel_line =  	16'b0011110011100000;
		12'h688:	pixel_line =  	16'b0011100001110000;
		12'h689:	pixel_line =  	16'b0011100000111000;
		12'h68A:	pixel_line =  	16'b0011100000111000;
		12'h68B:	pixel_line =  	16'b0011100000111000;
		12'h68C:	pixel_line =  	16'b0011100000111000;
		12'h68D:	pixel_line =  	16'b0000000000000000;
		12'h68E:	pixel_line =  	16'b0000000000000000;
		12'h68F:	pixel_line =  	16'b0000000000000000;

		12'h690:	pixel_line =  	16'b0000111100000000;  // i in ASCII
		12'h691:	pixel_line =  	16'b0000111100000000;
		12'h692:	pixel_line =  	16'b0000000000000000;
		12'h693:	pixel_line =  	16'b0000000000000000;
		12'h694:	pixel_line =  	16'b0011111100000000;
		12'h695:	pixel_line =  	16'b0011111100000000;
		12'h696:	pixel_line =  	16'b0000111100000000;
		12'h697:	pixel_line =  	16'b0000111100000000;
		12'h698:	pixel_line =  	16'b0000111100000000;
		12'h699:	pixel_line =  	16'b0000111100000000;
		12'h69A:	pixel_line =  	16'b0000111100000000;
		12'h69B:	pixel_line =  	16'b0011111111100000;
		12'h69C:	pixel_line =  	16'b0011111111100000;
		12'h69D:	pixel_line =  	16'b0000000000000000;
		12'h69E:	pixel_line =  	16'b0000000000000000;
		12'h69F:	pixel_line =  	16'b0000000000000000;

		12'h6A0:	pixel_line =  	16'b0000000001111000;  // j in ASCII
		12'h6A1:	pixel_line =  	16'b0000000001111000;
		12'h6A2:	pixel_line =  	16'b0000000000000000;
		12'h6A3:	pixel_line =  	16'b0000000000000000;
		12'h6A4:	pixel_line =  	16'b0001111111111000;
		12'h6A5:	pixel_line =  	16'b0001111111111000;
		12'h6A6:	pixel_line =  	16'b0000000000111000;
		12'h6A7:	pixel_line =  	16'b0000000000111000;
		12'h6A8:	pixel_line =  	16'b0000000000111000;
		12'h6A9:	pixel_line =  	16'b0000000000111000;
		12'h6AA:	pixel_line =  	16'b0000000000111000;
		12'h6AB:	pixel_line =  	16'b0011100001111000;
		12'h6AC:	pixel_line =  	16'b0011100011110000;
		12'h6AD:	pixel_line =  	16'b0001111111100000;
		12'h6AE:	pixel_line =  	16'b0000111111000000;
		12'h6AF:	pixel_line =  	16'b0000000000000000;

		12'h6B0:	pixel_line =  	16'b0000000000000000;  // k in ASCII 
		12'h6B1:	pixel_line =  	16'b0011100000000000;
		12'h6B2:	pixel_line =  	16'b0011100001110000;
		12'h6B3:	pixel_line =  	16'b0011100011100000;
		12'h6B4:	pixel_line =  	16'b0011100111000000;
		12'h6B5:	pixel_line =  	16'b0011101110000000;
		12'h6B6:	pixel_line =  	16'b0011111100000000;
		12'h6B7:	pixel_line =  	16'b0011111100000000;
		12'h6B8:	pixel_line =  	16'b0011101110000000;
		12'h6B9:	pixel_line =  	16'b0011100111000000;
		12'h6BA:	pixel_line =  	16'b0011100011100000;
		12'h6BB:	pixel_line =  	16'b0011100001110000;
		12'h6BC:	pixel_line =  	16'b0011100000111000;
		12'h6BD:	pixel_line =  	16'b0000000000000000;
		12'h6BE:	pixel_line =  	16'b0000000000000000;
		12'h6BF:	pixel_line =  	16'b0000000000000000;

		12'h6C0:	pixel_line =  	16'b0000000000000000;  // l in ASCII
		12'h6C1:	pixel_line =  	16'b0011111000000000;
		12'h6C2:	pixel_line =  	16'b0011111000000000;
		12'h6C3:	pixel_line =  	16'b0000111000000000;
		12'h6C4:	pixel_line =  	16'b0000111000000000;
		12'h6C5:	pixel_line =  	16'b0000111000000000;
		12'h6C6:	pixel_line =  	16'b0000111000000000;
		12'h6C7:	pixel_line =  	16'b0000111000000000;
		12'h6C8:	pixel_line =  	16'b0000111000000000;
		12'h6C9:	pixel_line =  	16'b0000111000000000;
		12'h6CA:	pixel_line =  	16'b0000111000000000;
		12'h6CB:	pixel_line =  	16'b0011111110000000;
		12'h6CC:	pixel_line =  	16'b0011111110000000;
		12'h6CD:	pixel_line =  	16'b0000000000000000;
		12'h6CE:	pixel_line =  	16'b0000000000000000;
		12'h6CF:	pixel_line =  	16'b0000000000000000;

		12'h6D0:	pixel_line =  	16'b0000000000000000;  // m in ASCII
		12'h6D1:	pixel_line =  	16'b0000000000000000;
		12'h6D2:	pixel_line =  	16'b0000000000000000;
		12'h6D3:	pixel_line =  	16'b0000000000000000;
		12'h6D4:	pixel_line =  	16'b0111110001110000;
		12'h6D5:	pixel_line =  	16'b0111111011111000;
		12'h6D6:	pixel_line =  	16'b0111001110011100;
		12'h6D7:	pixel_line =  	16'b0111001110011100;
		12'h6D8:	pixel_line =  	16'b0111001110011100;
		12'h6D9:	pixel_line =  	16'b0111001110011100;
		12'h6DA:	pixel_line =  	16'b0111001110011100;
		12'h6DB:	pixel_line =  	16'b0111001110011100;
		12'h6DC:	pixel_line =  	16'b0111001110011100;
		12'h6DD:	pixel_line =  	16'b0000000000000000;
		12'h6DE:	pixel_line =  	16'b0000000000000000;
		12'h6DF:	pixel_line =  	16'b0000000000000000;

		12'h6E0:	pixel_line =  	16'b0000000000000000;  // n in ASCII
		12'h6E1:	pixel_line =  	16'b0000000000000000;
		12'h6E2:	pixel_line =  	16'b0000000000000000;
		12'h6E3:	pixel_line =  	16'b0000000000000000;
		12'h6E4:	pixel_line =  	16'b0011100110000000;
		12'h6E5:	pixel_line =  	16'b0011101111100000;
		12'h6E6:	pixel_line =  	16'b0011111111110000;
		12'h6E7:	pixel_line =  	16'b0011110001111000;
		12'h6E8:	pixel_line =  	16'b0011100000111000;
		12'h6E9:	pixel_line =  	16'b0011100000011100;
		12'h6EA:	pixel_line =  	16'b0011100000011100;
		12'h6EB:	pixel_line =  	16'b0011100000011100;
		12'h6EC:	pixel_line =  	16'b0011100000011100;
		12'h6ED:	pixel_line =  	16'b0000000000000000;
		12'h6EE:	pixel_line =  	16'b0000000000000000;
		12'h6EF:	pixel_line =  	16'b0000000000000000;

		12'h6F0:	pixel_line =  	16'b0000000000000000;  // o in ASCII
		12'h6F1:	pixel_line =  	16'b0000000000000000;
		12'h6F2:	pixel_line =  	16'b0000000000000000;
		12'h6F3:	pixel_line =  	16'b0000011111100000;
		12'h6F4:	pixel_line =  	16'b0001111111111000;
		12'h6F5:	pixel_line =  	16'b0011110000111100;
		12'h6F6:	pixel_line =  	16'b0111100000011110;
		12'h6F7:	pixel_line =  	16'b0111000000001110;
		12'h6F8:	pixel_line =  	16'b0111000000001110;
		12'h6F9:	pixel_line =  	16'b0111100000011110;
		12'h6FA:	pixel_line =  	16'b0011110000111100;
		12'h6FB:	pixel_line =  	16'b0001111111111000;
		12'h6FC:	pixel_line =  	16'b0000111111110000;
		12'h6FD:	pixel_line =  	16'b0000000000000000;
		12'h6FE:	pixel_line =  	16'b0000000000000000;
		12'h6FF:	pixel_line =  	16'b0000000000000000;

		12'h700:	pixel_line =  	16'b0000000000000000;  // p in ASCII
		12'h701:	pixel_line =  	16'b0000000000000000;
		12'h702:	pixel_line =  	16'b0000000000000000;
		12'h703:	pixel_line =  	16'b0011100111000000;
		12'h704:	pixel_line =  	16'b0011101111110000;
		12'h705:	pixel_line =  	16'b0011111111111000;
		12'h706:	pixel_line =  	16'b0011110000111100;
		12'h707:	pixel_line =  	16'b0011100000011100;
		12'h708:	pixel_line =  	16'b0011100000111100;
		12'h709:	pixel_line =  	16'b0011100001111000;
		12'h70A:	pixel_line =  	16'b0011111111110000;
		12'h70B:	pixel_line =  	16'b0011110000000000;
		12'h70C:	pixel_line =  	16'b0011100000000000;
		12'h70D:	pixel_line =  	16'b0011100000000000;
		12'h70E:	pixel_line =  	16'b0011100000000000;
		12'h70F:	pixel_line =  	16'b0000000000000000;
		
		12'h710:	pixel_line =  	16'b0000000000000000;  // q in ASCII
		12'h711:	pixel_line =  	16'b0000000000000000;
		12'h712:	pixel_line =  	16'b0000000000000000;
		12'h713:	pixel_line =  	16'b0000011111111000;
		12'h714:	pixel_line =  	16'b0000111111111100;
		12'h715:	pixel_line =  	16'b0011110000111100;
		12'h716:	pixel_line =  	16'b0011100000011100;
		12'h717:	pixel_line =  	16'b0011100000011100;
		12'h718:	pixel_line =  	16'b0001110000111100;
		12'h719:	pixel_line =  	16'b0000111111111100;
		12'h71A:	pixel_line =  	16'b0000001111011100;
		12'h71B:	pixel_line =  	16'b0000000000011100;
		12'h71C:	pixel_line =  	16'b0000000000011100;
		12'h71D:	pixel_line =  	16'b0000000000011100;
		12'h71E:	pixel_line =  	16'b0000000000011100;
		12'h71F:	pixel_line =  	16'b0000000000000000;

		12'h720:	pixel_line =  	16'b0000000000000000;  // r in ASCII 
		12'h721:	pixel_line =  	16'b0000000000000000;
		12'h722:	pixel_line =  	16'b0000000000000000;
		12'h723:	pixel_line =  	16'b0011100110000000;
		12'h724:	pixel_line =  	16'b0011101111100000;
		12'h725:	pixel_line =  	16'b0011111111110000;
		12'h726:	pixel_line =  	16'b0011110001111000;
		12'h727:	pixel_line =  	16'b0011100000111000;
		12'h728:	pixel_line =  	16'b0011100000111000;
		12'h729:	pixel_line =  	16'b0011100000000000;
		12'h72A:	pixel_line =  	16'b0011100000000000;
		12'h72B:	pixel_line =  	16'b0011100000000000;
		12'h72C:	pixel_line =  	16'b0011100000000000;
		12'h72D:	pixel_line =  	16'b0000000000000000;
		12'h72E:	pixel_line =  	16'b0000000000000000;
		12'h72F:	pixel_line =  	16'b0000000000000000;

		12'h730:	pixel_line =  	16'b0000000000000000;  // s in ASCII
		12'h731:	pixel_line =  	16'b0000000000000000;
		12'h732:	pixel_line =  	16'b0000000000000000;
		12'h733:	pixel_line =  	16'b0000111111000000;
		12'h734:	pixel_line =  	16'b0011111111110000;
		12'h735:	pixel_line =  	16'b0111100000111000;
		12'h736:	pixel_line =  	16'b0011110000000000;
		12'h737:	pixel_line =  	16'b0000111100000000;
		12'h738:	pixel_line =  	16'b0000001111000000;
		12'h739:	pixel_line =  	16'b0000000111111000;
		12'h73A:	pixel_line =  	16'b0111000001111100;
		12'h73B:	pixel_line =  	16'b0011111111110000;
		12'h73C:	pixel_line =  	16'b0000111111000000;
		12'h73D:	pixel_line =  	16'b0000000000000000;
		12'h73E:	pixel_line =  	16'b0000000000000000;
		12'h73F:	pixel_line =  	16'b0000000000000000;

		12'h740:	pixel_line =  	16'b0000000000000000;  // t in ASCII
		12'h741:	pixel_line =  	16'b0000011100000000;
		12'h742:	pixel_line =  	16'b0000011100000000;
		12'h743:	pixel_line =  	16'b0001111111110000;
		12'h744:	pixel_line =  	16'b0001111111110000;
		12'h745:	pixel_line =  	16'b0000011100000000;
		12'h746:	pixel_line =  	16'b0000011100000000;
		12'h747:	pixel_line =  	16'b0000011100000000;
		12'h748:	pixel_line =  	16'b0000011100000000;
		12'h749:	pixel_line =  	16'b0000011100000000;
		12'h74A:	pixel_line =  	16'b0000011100000000;
		12'h74B:	pixel_line =  	16'b0000011111110000;
		12'h74C:	pixel_line =  	16'b0000001111110000;
		12'h74D:	pixel_line =  	16'b0000000000000000;
		12'h74E:	pixel_line =  	16'b0000000000000000;
		12'h74F:	pixel_line =  	16'b0000000000000000;

		12'h750:	pixel_line =  	16'b0000000000000000;  // u in ASCII
		12'h751:	pixel_line =  	16'b0000000000000000;
		12'h752:	pixel_line =  	16'b0000000000000000;
		12'h753:	pixel_line =  	16'b1111000011110000;
		12'h754:	pixel_line =  	16'b1111000011110000;
		12'h755:	pixel_line =  	16'b1111000011110000;
		12'h756:	pixel_line =  	16'b1111000011110000;
		12'h757:	pixel_line =  	16'b1111000011110000;
		12'h758:	pixel_line =  	16'b1111000011110000;
		12'h759:	pixel_line =  	16'b1111000011110000;
		12'h75A:	pixel_line =  	16'b1111100111111000;
		12'h75B:	pixel_line =  	16'b0111111101111100;
		12'h75C:	pixel_line =  	16'b0011111100111100;
		12'h75D:	pixel_line =  	16'b0000000000000000;
		12'h75E:	pixel_line =  	16'b0000000000000000;
		12'h75F:	pixel_line =  	16'b0000000000000000;

		12'h760:	pixel_line =  	16'b0000000000000000;  // v in ASCII
		12'h761:	pixel_line =  	16'b0000000000000000;
		12'h762:	pixel_line =  	16'b0000000000000000;
		12'h763:	pixel_line =  	16'b0000000000000000;
		12'h764:	pixel_line =  	16'b1110000000001110;
		12'h765:	pixel_line =  	16'b0111000000011100;
		12'h766:	pixel_line =  	16'b0111000000011100;
		12'h767:	pixel_line =  	16'b0011100000111000;
		12'h768:	pixel_line =  	16'b0011100000111000;
		12'h769:	pixel_line =  	16'b0001110001110000;
		12'h76A:	pixel_line =  	16'b0000110001100000;
		12'h76B:	pixel_line =  	16'b0000111011100000;
		12'h76C:	pixel_line =  	16'b0000011111000000;
		12'h76D:	pixel_line =  	16'b0000000000000000;
		12'h76E:	pixel_line =  	16'b0000000000000000;
		12'h76F:	pixel_line =  	16'b0000000000000000;

		12'h770:	pixel_line =  	16'b0000000000000000;  // w in ASCII 
		12'h771:	pixel_line =  	16'b0000000000000000;
		12'h772:	pixel_line =  	16'b0000000000000000;
		12'h773:	pixel_line =  	16'b0000000000000000;
		12'h774:	pixel_line =  	16'b0100000000000010;
		12'h775:	pixel_line =  	16'b0110000000000110;
		12'h776:	pixel_line =  	16'b0011000000001100;
		12'h777:	pixel_line =  	16'b0011100110011100;
		12'h778:	pixel_line =  	16'b0011101110111000;
		12'h779:	pixel_line =  	16'b0001111111110000;
		12'h77A:	pixel_line =  	16'b0000111011100000;
		12'h77B:	pixel_line =  	16'b0000110001100000;
		12'h77C:	pixel_line =  	16'b0000110001100000;
		12'h77D:	pixel_line =  	16'b0000000000000000;
		12'h77E:	pixel_line =  	16'b0000000000000000;
		12'h77F:	pixel_line =  	16'b0000000000000000;

		12'h780:	pixel_line =  	16'b0000000000000000;  // x in ASCII
		12'h781:	pixel_line =  	16'b0000000000000000;
		12'h782:	pixel_line =  	16'b0000000000000000;
		12'h783:	pixel_line =  	16'b0111000000011100;
		12'h784:	pixel_line =  	16'b0011100000111000;
		12'h785:	pixel_line =  	16'b0001110001110000;
		12'h786:	pixel_line =  	16'b0000111011100000;
		12'h787:	pixel_line =  	16'b0000011111000000;
		12'h788:	pixel_line =  	16'b0000011111000000;
		12'h789:	pixel_line =  	16'b0000111011100000;
		12'h78A:	pixel_line =  	16'b0001110001110000;
		12'h78B:	pixel_line =  	16'b0011100000111000;
		12'h78C:	pixel_line =  	16'b0111000000011100;
		12'h78D:	pixel_line =  	16'b0000000000000000;
		12'h78E:	pixel_line =  	16'b0000000000000000;
		12'h78F:	pixel_line =  	16'b0000000000000000;

		12'h790:	pixel_line =  	16'b0000000000000000;  // y in ASCII
		12'h791:	pixel_line =  	16'b0000000000000000;
		12'h792:	pixel_line =  	16'b0000000000000000;
		12'h793:	pixel_line =  	16'b0011100000001110;
		12'h794:	pixel_line =  	16'b0001110000011100;
		12'h795:	pixel_line =  	16'b0000111000111000;
		12'h796:	pixel_line =  	16'b0000011101110000;
		12'h797:	pixel_line =  	16'b0000001111100000;
		12'h798:	pixel_line =  	16'b0000000111100000;
		12'h799:	pixel_line =  	16'b0000001111000000;
		12'h79A:	pixel_line =  	16'b0000001110000000;
		12'h79B:	pixel_line =  	16'b0000111100000000;
		12'h79C:	pixel_line =  	16'b0011111000000000;
		12'h79D:	pixel_line =  	16'b0111100000000000;
		12'h79E:	pixel_line =  	16'b0000000000000000;
		12'h79F:	pixel_line =  	16'b0000000000000000;

		12'h7A0:	pixel_line =  	16'b0000000000000000;  // z in ASCII
		12'h7A1:	pixel_line =  	16'b0000000000000000;
		12'h7A2:	pixel_line =  	16'b0000000000000000;
		12'h7A3:	pixel_line =  	16'b1111111111110000;
		12'h7A4:	pixel_line =  	16'b1111111111110000;
		12'h7A5:	pixel_line =  	16'b1100001111100000;
		12'h7A6:	pixel_line =  	16'b1100011111000000;
		12'h7A7:	pixel_line =  	16'b0000111110000000;
		12'h7A8:	pixel_line =  	16'b0001111100000000;
		12'h7A9:	pixel_line =  	16'b0011111000110000;
		12'h7AA:	pixel_line =  	16'b0111110000110000;
		12'h7AB:	pixel_line =  	16'b1111111111110000;
		12'h7AC:	pixel_line =  	16'b1111111111110000;
		12'h7AD:	pixel_line =  	16'b0000000000000000;
		12'h7AE:	pixel_line =  	16'b0000000000000000;
		12'h7AF:	pixel_line =  	16'b0000000000000000;

		// empty
		default: pixel_line =  	16'b0000000000000000;

	endcase

  end








endmodule
